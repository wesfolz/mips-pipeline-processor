`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// ECE369 - Computer Architecture
// Module - data_memory.v
// Description - 32-Bit wide data memory. An example that shows how to prepare/initialize
// data memory
//
// INPUTS:-
// Address: 32-Bit address input port.
// WriteData: 32-Bit input port.
// Clk: 1-Bit Input clock signal.
// MemWrite: 1-Bit control signal for memory write.
// MemRead: 1-Bit control signal for memory read.
//
// OUTPUTS:-
// ReadData: 32-Bit registered output port.
//
// FUNCTIONALITY:-
// Design the above memory similar to the 'RegisterFile' model in the previous 
// assignment.  Create a memory and initialize it by reading from a test data.  
// The 'WriteData' value is written into the address 
// in the positive clock edge if 'MemWrite' 
// signal is 1. 'ReadData' is the value of memory location if 
// 'MemRead' is 1, otherwise, it is 0x00000000. The reading of memory is not 
// clocked.
////////////////////////////////////////////////////////////////////////////////

module DataMemory(Address, MemRead, ReadData); 

    input [31:0] Address;   // Input Address 
  //  input [31:0] WriteData; // Data that needs to be written into the address 
 //   input Clk;
 //   input MemWrite;         // Control signal for memory write 
    input MemRead;          // Control signal for memory read 
	// integer i;			
	

    output reg[31:0] ReadData; // Contents of memory location at Address

    reg [31:0] memory[0:1043];    // size needs to be adjusted based on the size of the test_data.txt
	
	 	 
	 initial begin
	 

		 

//result should be 28, 28
memory[0] = 32'h20;
memory[1] = 32'h20;
memory[2] = 32'h4;
memory[3] = 32'h4;
memory[4] = 32'h1;
memory[5] = 32'h1;
memory[6] = 32'h1;
memory[7] = 32'h1;
memory[8] = 32'h1;
memory[9] = 32'h1;
memory[10] = 32'h1;
memory[11] = 32'h1;
memory[12] = 32'h1;
memory[13] = 32'h1;
memory[14] = 32'h1;
memory[15] = 32'h1;
memory[16] = 32'h1;
memory[17] = 32'h1;
memory[18] = 32'h1;
memory[19] = 32'h1;
memory[20] = 32'h1;
memory[21] = 32'h1;
memory[22] = 32'h1;
memory[23] = 32'h1;
memory[24] = 32'h1;
memory[25] = 32'h1;
memory[26] = 32'h1;
memory[27] = 32'h1;
memory[28] = 32'h1;
memory[29] = 32'h1;
memory[30] = 32'h1;
memory[31] = 32'h1;
memory[32] = 32'h1;
memory[33] = 32'h1;
memory[34] = 32'h1;
memory[35] = 32'h1;
memory[36] = 32'h1;
memory[37] = 32'h1;
memory[38] = 32'h1;
memory[39] = 32'h1;
memory[40] = 32'h1;
memory[41] = 32'h1;
memory[42] = 32'h1;
memory[43] = 32'h1;
memory[44] = 32'h1;
memory[45] = 32'h1;
memory[46] = 32'h1;
memory[47] = 32'h1;
memory[48] = 32'h1;
memory[49] = 32'h1;
memory[50] = 32'h1;
memory[51] = 32'h1;
memory[52] = 32'h1;
memory[53] = 32'h1;
memory[54] = 32'h1;
memory[55] = 32'h1;
memory[56] = 32'h1;
memory[57] = 32'h1;
memory[58] = 32'h1;
memory[59] = 32'h1;
memory[60] = 32'h1;
memory[61] = 32'h1;
memory[62] = 32'h1;
memory[63] = 32'h1;
memory[64] = 32'h1;
memory[65] = 32'h1;
memory[66] = 32'h1;
memory[67] = 32'h1;
memory[68] = 32'h1;
memory[69] = 32'h1;
memory[70] = 32'h1;
memory[71] = 32'h1;
memory[72] = 32'h1;
memory[73] = 32'h1;
memory[74] = 32'h1;
memory[75] = 32'h1;
memory[76] = 32'h1;
memory[77] = 32'h1;
memory[78] = 32'h1;
memory[79] = 32'h1;
memory[80] = 32'h1;
memory[81] = 32'h1;
memory[82] = 32'h1;
memory[83] = 32'h1;
memory[84] = 32'h1;
memory[85] = 32'h1;
memory[86] = 32'h1;
memory[87] = 32'h1;
memory[88] = 32'h1;
memory[89] = 32'h1;
memory[90] = 32'h1;
memory[91] = 32'h1;
memory[92] = 32'h1;
memory[93] = 32'h1;
memory[94] = 32'h1;
memory[95] = 32'h1;
memory[96] = 32'h1;
memory[97] = 32'h1;
memory[98] = 32'h1;
memory[99] = 32'h1;
memory[100] = 32'h1;
memory[101] = 32'h1;
memory[102] = 32'h1;
memory[103] = 32'h1;
memory[104] = 32'h1;
memory[105] = 32'h1;
memory[106] = 32'h1;
memory[107] = 32'h1;
memory[108] = 32'h1;
memory[109] = 32'h1;
memory[110] = 32'h1;
memory[111] = 32'h1;
memory[112] = 32'h1;
memory[113] = 32'h1;
memory[114] = 32'h1;
memory[115] = 32'h1;
memory[116] = 32'h1;
memory[117] = 32'h1;
memory[118] = 32'h1;
memory[119] = 32'h1;
memory[120] = 32'h1;
memory[121] = 32'h1;
memory[122] = 32'h1;
memory[123] = 32'h1;
memory[124] = 32'h1;
memory[125] = 32'h1;
memory[126] = 32'h1;
memory[127] = 32'h1;
memory[128] = 32'h1;
memory[129] = 32'h1;
memory[130] = 32'h1;
memory[131] = 32'h1;
memory[132] = 32'h1;
memory[133] = 32'h1;
memory[134] = 32'h1;
memory[135] = 32'h1;
memory[136] = 32'h1;
memory[137] = 32'h1;
memory[138] = 32'h1;
memory[139] = 32'h1;
memory[140] = 32'h1;
memory[141] = 32'h1;
memory[142] = 32'h1;
memory[143] = 32'h1;
memory[144] = 32'h1;
memory[145] = 32'h1;
memory[146] = 32'h1;
memory[147] = 32'h1;
memory[148] = 32'h1;
memory[149] = 32'h1;
memory[150] = 32'h1;
memory[151] = 32'h1;
memory[152] = 32'h1;
memory[153] = 32'h1;
memory[154] = 32'h1;
memory[155] = 32'h1;
memory[156] = 32'h1;
memory[157] = 32'h1;
memory[158] = 32'h1;
memory[159] = 32'h1;
memory[160] = 32'h1;
memory[161] = 32'h1;
memory[162] = 32'h1;
memory[163] = 32'h1;
memory[164] = 32'h1;
memory[165] = 32'h1;
memory[166] = 32'h1;
memory[167] = 32'h1;
memory[168] = 32'h1;
memory[169] = 32'h1;
memory[170] = 32'h1;
memory[171] = 32'h1;
memory[172] = 32'h1;
memory[173] = 32'h1;
memory[174] = 32'h1;
memory[175] = 32'h1;
memory[176] = 32'h1;
memory[177] = 32'h1;
memory[178] = 32'h1;
memory[179] = 32'h1;
memory[180] = 32'h1;
memory[181] = 32'h1;
memory[182] = 32'h1;
memory[183] = 32'h1;
memory[184] = 32'hb;
memory[185] = 32'hb;
memory[186] = 32'hb;
memory[187] = 32'hb;
memory[188] = 32'hb;
memory[189] = 32'hb;
memory[190] = 32'hb;
memory[191] = 32'hb;
memory[192] = 32'hb;
memory[193] = 32'hb;
memory[194] = 32'hb;
memory[195] = 32'hb;
memory[196] = 32'h1;
memory[197] = 32'h1;
memory[198] = 32'h1;
memory[199] = 32'h1;
memory[200] = 32'h1;
memory[201] = 32'h1;
memory[202] = 32'h1;
memory[203] = 32'h1;
memory[204] = 32'h1;
memory[205] = 32'h1;
memory[206] = 32'h1;
memory[207] = 32'h1;
memory[208] = 32'h1;
memory[209] = 32'h1;
memory[210] = 32'h1;
memory[211] = 32'h1;
memory[212] = 32'h1;
memory[213] = 32'h1;
memory[214] = 32'h1;
memory[215] = 32'h1;
memory[216] = 32'hb;
memory[217] = 32'hb;
memory[218] = 32'hb;
memory[219] = 32'hb;
memory[220] = 32'hb;
memory[221] = 32'hb;
memory[222] = 32'hb;
memory[223] = 32'hb;
memory[224] = 32'hb;
memory[225] = 32'hb;
memory[226] = 32'hb;
memory[227] = 32'hb;
memory[228] = 32'h1;
memory[229] = 32'h1;
memory[230] = 32'h1;
memory[231] = 32'h1;
memory[232] = 32'h1;
memory[233] = 32'h1;
memory[234] = 32'h1;
memory[235] = 32'h1;
memory[236] = 32'h1;
memory[237] = 32'h1;
memory[238] = 32'h1;
memory[239] = 32'h1;
memory[240] = 32'h1;
memory[241] = 32'h1;
memory[242] = 32'h1;
memory[243] = 32'h1;
memory[244] = 32'h1;
memory[245] = 32'h1;
memory[246] = 32'h1;
memory[247] = 32'h1;
memory[248] = 32'hb;
memory[249] = 32'hb;
memory[250] = 32'hb;
memory[251] = 32'hb;
memory[252] = 32'hb;
memory[253] = 32'hb;
memory[254] = 32'hb;
memory[255] = 32'hb;
memory[256] = 32'hb;
memory[257] = 32'hb;
memory[258] = 32'hb;
memory[259] = 32'hb;
memory[260] = 32'h1;
memory[261] = 32'h1;
memory[262] = 32'h1;
memory[263] = 32'h1;
memory[264] = 32'h1;
memory[265] = 32'h1;
memory[266] = 32'h1;
memory[267] = 32'h1;
memory[268] = 32'h1;
memory[269] = 32'h1;
memory[270] = 32'h1;
memory[271] = 32'h1;
memory[272] = 32'h1;
memory[273] = 32'h1;
memory[274] = 32'h1;
memory[275] = 32'h1;
memory[276] = 32'h1;
memory[277] = 32'h1;
memory[278] = 32'h1;
memory[279] = 32'h1;
memory[280] = 32'hb;
memory[281] = 32'hb;
memory[282] = 32'hb;
memory[283] = 32'hb;
memory[284] = 32'hb;
memory[285] = 32'hb;
memory[286] = 32'hb;
memory[287] = 32'hb;
memory[288] = 32'hb;
memory[289] = 32'hb;
memory[290] = 32'hb;
memory[291] = 32'hb;
memory[292] = 32'h1;
memory[293] = 32'h1;
memory[294] = 32'h1;
memory[295] = 32'h1;
memory[296] = 32'h1;
memory[297] = 32'h1;
memory[298] = 32'h1;
memory[299] = 32'h1;
memory[300] = 32'h1;
memory[301] = 32'h1;
memory[302] = 32'h1;
memory[303] = 32'h1;
memory[304] = 32'h1;
memory[305] = 32'h1;
memory[306] = 32'h1;
memory[307] = 32'h1;
memory[308] = 32'h1;
memory[309] = 32'h1;
memory[310] = 32'h1;
memory[311] = 32'h1;
memory[312] = 32'hb;
memory[313] = 32'hb;
memory[314] = 32'hb;
memory[315] = 32'hb;
memory[316] = 32'hb;
memory[317] = 32'hb;
memory[318] = 32'hb;
memory[319] = 32'hb;
memory[320] = 32'hb;
memory[321] = 32'hb;
memory[322] = 32'hb;
memory[323] = 32'hb;
memory[324] = 32'h1;
memory[325] = 32'h1;
memory[326] = 32'h1;
memory[327] = 32'h1;
memory[328] = 32'h1;
memory[329] = 32'h1;
memory[330] = 32'h1;
memory[331] = 32'h1;
memory[332] = 32'h1;
memory[333] = 32'h1;
memory[334] = 32'h1;
memory[335] = 32'h1;
memory[336] = 32'h1;
memory[337] = 32'h1;
memory[338] = 32'h1;
memory[339] = 32'h1;
memory[340] = 32'h1;
memory[341] = 32'h1;
memory[342] = 32'h1;
memory[343] = 32'h1;
memory[344] = 32'hb;
memory[345] = 32'hb;
memory[346] = 32'hb;
memory[347] = 32'hb;
memory[348] = 32'hb;
memory[349] = 32'hb;
memory[350] = 32'hb;
memory[351] = 32'hb;
memory[352] = 32'hb;
memory[353] = 32'hb;
memory[354] = 32'hb;
memory[355] = 32'hb;
memory[356] = 32'h1;
memory[357] = 32'h1;
memory[358] = 32'h1;
memory[359] = 32'h1;
memory[360] = 32'h1;
memory[361] = 32'h1;
memory[362] = 32'h1;
memory[363] = 32'h1;
memory[364] = 32'h1;
memory[365] = 32'h1;
memory[366] = 32'h1;
memory[367] = 32'h1;
memory[368] = 32'h1;
memory[369] = 32'h1;
memory[370] = 32'h1;
memory[371] = 32'h1;
memory[372] = 32'h1;
memory[373] = 32'h1;
memory[374] = 32'h1;
memory[375] = 32'h1;
memory[376] = 32'hb;
memory[377] = 32'hb;
memory[378] = 32'hb;
memory[379] = 32'hb;
memory[380] = 32'hb;
memory[381] = 32'hb;
memory[382] = 32'hb;
memory[383] = 32'hb;
memory[384] = 32'hb;
memory[385] = 32'hb;
memory[386] = 32'hb;
memory[387] = 32'hb;
memory[388] = 32'h1;
memory[389] = 32'h1;
memory[390] = 32'h1;
memory[391] = 32'h1;
memory[392] = 32'h1;
memory[393] = 32'h1;
memory[394] = 32'h1;
memory[395] = 32'h1;
memory[396] = 32'h1;
memory[397] = 32'h1;
memory[398] = 32'h1;
memory[399] = 32'h1;
memory[400] = 32'h1;
memory[401] = 32'h1;
memory[402] = 32'h1;
memory[403] = 32'h1;
memory[404] = 32'h1;
memory[405] = 32'h1;
memory[406] = 32'h1;
memory[407] = 32'h1;
memory[408] = 32'hb;
memory[409] = 32'hb;
memory[410] = 32'hb;
memory[411] = 32'hb;
memory[412] = 32'hb;
memory[413] = 32'hb;
memory[414] = 32'hb;
memory[415] = 32'hb;
memory[416] = 32'hb;
memory[417] = 32'hb;
memory[418] = 32'hb;
memory[419] = 32'hb;
memory[420] = 32'h1;
memory[421] = 32'h1;
memory[422] = 32'h1;
memory[423] = 32'h1;
memory[424] = 32'h1;
memory[425] = 32'h1;
memory[426] = 32'h1;
memory[427] = 32'h1;
memory[428] = 32'h1;
memory[429] = 32'h1;
memory[430] = 32'h1;
memory[431] = 32'h1;
memory[432] = 32'h1;
memory[433] = 32'h1;
memory[434] = 32'h1;
memory[435] = 32'h1;
memory[436] = 32'h1;
memory[437] = 32'h1;
memory[438] = 32'h1;
memory[439] = 32'h1;
memory[440] = 32'hb;
memory[441] = 32'hb;
memory[442] = 32'hb;
memory[443] = 32'hb;
memory[444] = 32'hb;
memory[445] = 32'hb;
memory[446] = 32'hb;
memory[447] = 32'hb;
memory[448] = 32'hb;
memory[449] = 32'hb;
memory[450] = 32'hb;
memory[451] = 32'hb;
memory[452] = 32'h1;
memory[453] = 32'h1;
memory[454] = 32'h1;
memory[455] = 32'h1;
memory[456] = 32'h1;
memory[457] = 32'h1;
memory[458] = 32'h1;
memory[459] = 32'h1;
memory[460] = 32'h1;
memory[461] = 32'h1;
memory[462] = 32'h1;
memory[463] = 32'h1;
memory[464] = 32'h1;
memory[465] = 32'h1;
memory[466] = 32'h1;
memory[467] = 32'h1;
memory[468] = 32'h1;
memory[469] = 32'h1;
memory[470] = 32'h1;
memory[471] = 32'h1;
memory[472] = 32'hb;
memory[473] = 32'hb;
memory[474] = 32'hb;
memory[475] = 32'hb;
memory[476] = 32'hb;
memory[477] = 32'hb;
memory[478] = 32'hb;
memory[479] = 32'hb;
memory[480] = 32'hb;
memory[481] = 32'hb;
memory[482] = 32'hb;
memory[483] = 32'hb;
memory[484] = 32'h1;
memory[485] = 32'h1;
memory[486] = 32'h1;
memory[487] = 32'h1;
memory[488] = 32'h1;
memory[489] = 32'h1;
memory[490] = 32'h1;
memory[491] = 32'h1;
memory[492] = 32'h1;
memory[493] = 32'h1;
memory[494] = 32'h1;
memory[495] = 32'h1;
memory[496] = 32'h1;
memory[497] = 32'h1;
memory[498] = 32'h1;
memory[499] = 32'h1;
memory[500] = 32'h1;
memory[501] = 32'h1;
memory[502] = 32'h1;
memory[503] = 32'h1;
memory[504] = 32'hb;
memory[505] = 32'hb;
memory[506] = 32'hb;
memory[507] = 32'hb;
memory[508] = 32'hb;
memory[509] = 32'hb;
memory[510] = 32'hb;
memory[511] = 32'hb;
memory[512] = 32'hb;
memory[513] = 32'hb;
memory[514] = 32'hb;
memory[515] = 32'hb;
memory[516] = 32'h1;
memory[517] = 32'h1;
memory[518] = 32'h1;
memory[519] = 32'h1;
memory[520] = 32'h1;
memory[521] = 32'h1;
memory[522] = 32'h1;
memory[523] = 32'h1;
memory[524] = 32'h1;
memory[525] = 32'h1;
memory[526] = 32'h1;
memory[527] = 32'h1;
memory[528] = 32'h1;
memory[529] = 32'h1;
memory[530] = 32'h1;
memory[531] = 32'h1;
memory[532] = 32'h1;
memory[533] = 32'h1;
memory[534] = 32'h1;
memory[535] = 32'h1;
memory[536] = 32'hb;
memory[537] = 32'hb;
memory[538] = 32'hb;
memory[539] = 32'hb;
memory[540] = 32'hb;
memory[541] = 32'hb;
memory[542] = 32'hb;
memory[543] = 32'hb;
memory[544] = 32'hb;
memory[545] = 32'hb;
memory[546] = 32'hb;
memory[547] = 32'hb;
memory[548] = 32'h1;
memory[549] = 32'h1;
memory[550] = 32'h1;
memory[551] = 32'h1;
memory[552] = 32'h1;
memory[553] = 32'h1;
memory[554] = 32'h1;
memory[555] = 32'h1;
memory[556] = 32'h1;
memory[557] = 32'h1;
memory[558] = 32'h1;
memory[559] = 32'h1;
memory[560] = 32'h1;
memory[561] = 32'h1;
memory[562] = 32'h1;
memory[563] = 32'h1;
memory[564] = 32'h1;
memory[565] = 32'h1;
memory[566] = 32'h1;
memory[567] = 32'h1;
memory[568] = 32'hb;
memory[569] = 32'hb;
memory[570] = 32'hb;
memory[571] = 32'hb;
memory[572] = 32'hb;
memory[573] = 32'hb;
memory[574] = 32'hb;
memory[575] = 32'hb;
memory[576] = 32'hb;
memory[577] = 32'hb;
memory[578] = 32'hb;
memory[579] = 32'hb;
memory[580] = 32'h1;
memory[581] = 32'h1;
memory[582] = 32'h1;
memory[583] = 32'h1;
memory[584] = 32'h1;
memory[585] = 32'h1;
memory[586] = 32'h1;
memory[587] = 32'h1;
memory[588] = 32'h1;
memory[589] = 32'h1;
memory[590] = 32'h1;
memory[591] = 32'h1;
memory[592] = 32'h1;
memory[593] = 32'h1;
memory[594] = 32'h1;
memory[595] = 32'h1;
memory[596] = 32'h1;
memory[597] = 32'h1;
memory[598] = 32'h1;
memory[599] = 32'h1;
memory[600] = 32'hb;
memory[601] = 32'hb;
memory[602] = 32'hb;
memory[603] = 32'hb;
memory[604] = 32'hb;
memory[605] = 32'hb;
memory[606] = 32'hb;
memory[607] = 32'hb;
memory[608] = 32'hb;
memory[609] = 32'hb;
memory[610] = 32'hb;
memory[611] = 32'hb;
memory[612] = 32'h1;
memory[613] = 32'h1;
memory[614] = 32'h1;
memory[615] = 32'h1;
memory[616] = 32'h1;
memory[617] = 32'h1;
memory[618] = 32'h1;
memory[619] = 32'h1;
memory[620] = 32'h1;
memory[621] = 32'h1;
memory[622] = 32'h1;
memory[623] = 32'h1;
memory[624] = 32'h1;
memory[625] = 32'h1;
memory[626] = 32'h1;
memory[627] = 32'h1;
memory[628] = 32'h1;
memory[629] = 32'h1;
memory[630] = 32'h1;
memory[631] = 32'h1;
memory[632] = 32'ha;
memory[633] = 32'ha;
memory[634] = 32'ha;
memory[635] = 32'ha;
memory[636] = 32'ha;
memory[637] = 32'ha;
memory[638] = 32'ha;
memory[639] = 32'ha;
memory[640] = 32'ha;
memory[641] = 32'ha;
memory[642] = 32'ha;
memory[643] = 32'ha;
memory[644] = 32'h1;
memory[645] = 32'h1;
memory[646] = 32'h1;
memory[647] = 32'h1;
memory[648] = 32'h1;
memory[649] = 32'h1;
memory[650] = 32'h1;
memory[651] = 32'h1;
memory[652] = 32'h1;
memory[653] = 32'h1;
memory[654] = 32'h1;
memory[655] = 32'h1;
memory[656] = 32'h1;
memory[657] = 32'h1;
memory[658] = 32'h1;
memory[659] = 32'h1;
memory[660] = 32'h1;
memory[661] = 32'h1;
memory[662] = 32'h1;
memory[663] = 32'h1;
memory[664] = 32'ha;
memory[665] = 32'ha;
memory[666] = 32'ha;
memory[667] = 32'ha;
memory[668] = 32'ha;
memory[669] = 32'ha;
memory[670] = 32'ha;
memory[671] = 32'ha;
memory[672] = 32'ha;
memory[673] = 32'ha;
memory[674] = 32'ha;
memory[675] = 32'ha;
memory[676] = 32'h1;
memory[677] = 32'h1;
memory[678] = 32'h1;
memory[679] = 32'h1;
memory[680] = 32'h1;
memory[681] = 32'h1;
memory[682] = 32'h1;
memory[683] = 32'h1;
memory[684] = 32'h1;
memory[685] = 32'h1;
memory[686] = 32'h1;
memory[687] = 32'h1;
memory[688] = 32'h1;
memory[689] = 32'h1;
memory[690] = 32'h1;
memory[691] = 32'h1;
memory[692] = 32'h1;
memory[693] = 32'h1;
memory[694] = 32'h1;
memory[695] = 32'h1;
memory[696] = 32'h1;
memory[697] = 32'h1;
memory[698] = 32'h1;
memory[699] = 32'h1;
memory[700] = 32'h1;
memory[701] = 32'h1;
memory[702] = 32'h1;
memory[703] = 32'h1;
memory[704] = 32'h1;
memory[705] = 32'h1;
memory[706] = 32'h1;
memory[707] = 32'h1;
memory[708] = 32'h1;
memory[709] = 32'h1;
memory[710] = 32'h1;
memory[711] = 32'h1;
memory[712] = 32'h1;
memory[713] = 32'h1;
memory[714] = 32'h1;
memory[715] = 32'h1;
memory[716] = 32'h1;
memory[717] = 32'h1;
memory[718] = 32'h1;
memory[719] = 32'h1;
memory[720] = 32'h1;
memory[721] = 32'h1;
memory[722] = 32'h1;
memory[723] = 32'h1;
memory[724] = 32'h1;
memory[725] = 32'h1;
memory[726] = 32'h1;
memory[727] = 32'h1;
memory[728] = 32'h1;
memory[729] = 32'h1;
memory[730] = 32'h1;
memory[731] = 32'h1;
memory[732] = 32'h1;
memory[733] = 32'h1;
memory[734] = 32'h1;
memory[735] = 32'h1;
memory[736] = 32'h1;
memory[737] = 32'h1;
memory[738] = 32'h1;
memory[739] = 32'h1;
memory[740] = 32'h1;
memory[741] = 32'h1;
memory[742] = 32'h1;
memory[743] = 32'h1;
memory[744] = 32'h1;
memory[745] = 32'h1;
memory[746] = 32'h1;
memory[747] = 32'h1;
memory[748] = 32'h1;
memory[749] = 32'h1;
memory[750] = 32'h1;
memory[751] = 32'h1;
memory[752] = 32'h1;
memory[753] = 32'h1;
memory[754] = 32'h1;
memory[755] = 32'h1;
memory[756] = 32'h1;
memory[757] = 32'h1;
memory[758] = 32'h1;
memory[759] = 32'h1;
memory[760] = 32'h1;
memory[761] = 32'h1;
memory[762] = 32'h1;
memory[763] = 32'h1;
memory[764] = 32'h1;
memory[765] = 32'h1;
memory[766] = 32'h1;
memory[767] = 32'h1;
memory[768] = 32'h1;
memory[769] = 32'h1;
memory[770] = 32'h1;
memory[771] = 32'h1;
memory[772] = 32'h1;
memory[773] = 32'h1;
memory[774] = 32'h1;
memory[775] = 32'h1;
memory[776] = 32'h1;
memory[777] = 32'h1;
memory[778] = 32'h1;
memory[779] = 32'h1;
memory[780] = 32'h1;
memory[781] = 32'h1;
memory[782] = 32'h1;
memory[783] = 32'h1;
memory[784] = 32'h1;
memory[785] = 32'h1;
memory[786] = 32'h1;
memory[787] = 32'h1;
memory[788] = 32'h1;
memory[789] = 32'h1;
memory[790] = 32'h1;
memory[791] = 32'h1;
memory[792] = 32'h1;
memory[793] = 32'h1;
memory[794] = 32'h1;
memory[795] = 32'h1;
memory[796] = 32'h1;
memory[797] = 32'h1;
memory[798] = 32'h1;
memory[799] = 32'h1;
memory[800] = 32'h1;
memory[801] = 32'h1;
memory[802] = 32'h1;
memory[803] = 32'h1;
memory[804] = 32'h1;
memory[805] = 32'h1;
memory[806] = 32'h1;
memory[807] = 32'h1;
memory[808] = 32'h1;
memory[809] = 32'h1;
memory[810] = 32'h1;
memory[811] = 32'h1;
memory[812] = 32'h1;
memory[813] = 32'h1;
memory[814] = 32'h1;
memory[815] = 32'h1;
memory[816] = 32'h1;
memory[817] = 32'h1;
memory[818] = 32'h1;
memory[819] = 32'h1;
memory[820] = 32'h1;
memory[821] = 32'h1;
memory[822] = 32'h1;
memory[823] = 32'h1;
memory[824] = 32'h1;
memory[825] = 32'h1;
memory[826] = 32'h1;
memory[827] = 32'h1;
memory[828] = 32'h1;
memory[829] = 32'h1;
memory[830] = 32'h1;
memory[831] = 32'h1;
memory[832] = 32'h1;
memory[833] = 32'h1;
memory[834] = 32'h1;
memory[835] = 32'h1;
memory[836] = 32'h1;
memory[837] = 32'h1;
memory[838] = 32'h1;
memory[839] = 32'h1;
memory[840] = 32'h1;
memory[841] = 32'h1;
memory[842] = 32'h1;
memory[843] = 32'h1;
memory[844] = 32'h1;
memory[845] = 32'h1;
memory[846] = 32'h1;
memory[847] = 32'h1;
memory[848] = 32'h1;
memory[849] = 32'h1;
memory[850] = 32'h1;
memory[851] = 32'h1;
memory[852] = 32'h1;
memory[853] = 32'h1;
memory[854] = 32'h1;
memory[855] = 32'h1;
memory[856] = 32'h1;
memory[857] = 32'h1;
memory[858] = 32'h1;
memory[859] = 32'h1;
memory[860] = 32'h1;
memory[861] = 32'h1;
memory[862] = 32'h1;
memory[863] = 32'h1;
memory[864] = 32'h1;
memory[865] = 32'h1;
memory[866] = 32'h1;
memory[867] = 32'h1;
memory[868] = 32'h1;
memory[869] = 32'h1;
memory[870] = 32'h1;
memory[871] = 32'h1;
memory[872] = 32'h1;
memory[873] = 32'h1;
memory[874] = 32'h1;
memory[875] = 32'h1;
memory[876] = 32'h1;
memory[877] = 32'h1;
memory[878] = 32'h1;
memory[879] = 32'h1;
memory[880] = 32'h1;
memory[881] = 32'h1;
memory[882] = 32'h1;
memory[883] = 32'h1;
memory[884] = 32'h1;
memory[885] = 32'h1;
memory[886] = 32'h1;
memory[887] = 32'h1;
memory[888] = 32'h1;
memory[889] = 32'h1;
memory[890] = 32'h1;
memory[891] = 32'h1;
memory[892] = 32'h1;
memory[893] = 32'h1;
memory[894] = 32'h1;
memory[895] = 32'h1;
memory[896] = 32'h1;
memory[897] = 32'h1;
memory[898] = 32'h1;
memory[899] = 32'h1;
memory[900] = 32'h1;
memory[901] = 32'h1;
memory[902] = 32'h1;
memory[903] = 32'h1;
memory[904] = 32'h1;
memory[905] = 32'h1;
memory[906] = 32'h1;
memory[907] = 32'h1;
memory[908] = 32'h1;
memory[909] = 32'h1;
memory[910] = 32'h1;
memory[911] = 32'h1;
memory[912] = 32'h1;
memory[913] = 32'h1;
memory[914] = 32'h1;
memory[915] = 32'h1;
memory[916] = 32'h1;
memory[917] = 32'h1;
memory[918] = 32'h1;
memory[919] = 32'h1;
memory[920] = 32'h1;
memory[921] = 32'h1;
memory[922] = 32'h1;
memory[923] = 32'h1;
memory[924] = 32'h1;
memory[925] = 32'h1;
memory[926] = 32'h1;
memory[927] = 32'h1;
memory[928] = 32'ha;
memory[929] = 32'ha;
memory[930] = 32'ha;
memory[931] = 32'ha;
memory[932] = 32'h1;
memory[933] = 32'h1;
memory[934] = 32'h1;
memory[935] = 32'h1;
memory[936] = 32'h1;
memory[937] = 32'h1;
memory[938] = 32'h1;
memory[939] = 32'h1;
memory[940] = 32'h1;
memory[941] = 32'h1;
memory[942] = 32'h1;
memory[943] = 32'h1;
memory[944] = 32'h1;
memory[945] = 32'h1;
memory[946] = 32'h1;
memory[947] = 32'h1;
memory[948] = 32'h1;
memory[949] = 32'h1;
memory[950] = 32'h1;
memory[951] = 32'h1;
memory[952] = 32'h1;
memory[953] = 32'h1;
memory[954] = 32'h1;
memory[955] = 32'h1;
memory[956] = 32'h1;
memory[957] = 32'h1;
memory[958] = 32'h1;
memory[959] = 32'h1;
memory[960] = 32'ha;
memory[961] = 32'ha;
memory[962] = 32'ha;
memory[963] = 32'ha;
memory[964] = 32'h1;
memory[965] = 32'h1;
memory[966] = 32'h1;
memory[967] = 32'h1;
memory[968] = 32'h1;
memory[969] = 32'h1;
memory[970] = 32'h1;
memory[971] = 32'h1;
memory[972] = 32'h1;
memory[973] = 32'h1;
memory[974] = 32'h1;
memory[975] = 32'h1;
memory[976] = 32'h1;
memory[977] = 32'h1;
memory[978] = 32'h1;
memory[979] = 32'h1;
memory[980] = 32'h1;
memory[981] = 32'h1;
memory[982] = 32'h1;
memory[983] = 32'h1;
memory[984] = 32'h1;
memory[985] = 32'h1;
memory[986] = 32'h1;
memory[987] = 32'h1;
memory[988] = 32'h1;
memory[989] = 32'h1;
memory[990] = 32'h1;
memory[991] = 32'h1;
memory[992] = 32'ha;
memory[993] = 32'ha;
memory[994] = 32'ha;
memory[995] = 32'ha;
memory[996] = 32'h1;
memory[997] = 32'h1;
memory[998] = 32'h1;
memory[999] = 32'h1;
memory[1000] = 32'h1;
memory[1001] = 32'h1;
memory[1002] = 32'h1;
memory[1003] = 32'h1;
memory[1004] = 32'h1;
memory[1005] = 32'h1;
memory[1006] = 32'h1;
memory[1007] = 32'h1;
memory[1008] = 32'h1;
memory[1009] = 32'h1;
memory[1010] = 32'h1;
memory[1011] = 32'h1;
memory[1012] = 32'h1;
memory[1013] = 32'h1;
memory[1014] = 32'h1;
memory[1015] = 32'h1;
memory[1016] = 32'h1;
memory[1017] = 32'h1;
memory[1018] = 32'h1;
memory[1019] = 32'h1;
memory[1020] = 32'h1;
memory[1021] = 32'h1;
memory[1022] = 32'h1;
memory[1023] = 32'h1;
memory[1024] = 32'ha;
memory[1025] = 32'ha;
memory[1026] = 32'ha;
memory[1027] = 32'ha;
memory[1028] = 32'ha;
memory[1029] = 32'ha;
memory[1030] = 32'ha;
memory[1031] = 32'ha;
memory[1032] = 32'ha;
memory[1033] = 32'ha;
memory[1034] = 32'ha;
memory[1035] = 32'ha;
memory[1036] = 32'ha;
memory[1037] = 32'ha;
memory[1038] = 32'ha;
memory[1039] = 32'ha;
memory[1040] = 32'ha;
memory[1041] = 32'ha;
memory[1042] = 32'ha;
memory[1043] = 32'ha;



		
	 
	 
	 /*
	 
	 
	 //TestCase for Branches, Jump, SW, LW 
	
			//Initialize your Datamemory first as the following:		
			memory[1] <= 32'h00000001;
			memory[2] <= 32'hffffffff;
		
			
			//memory[*] <= 0, where * represents all the other indexes other than 1 and 2
			memory[0] <= 0;
			for(i=3;i<=31;i=i+1)begin			
				memory[i] <= 0;
			end
			
	 //End of TestCase for Branches, Jump, SW, LW
	 */
	
	 end 
	 /*
    always @(posedge Clk) begin      //memory write
        if (MemWrite==1)
            memory[Address[31:2]] <= WriteData;
    end
*/

    always @(Address or MemRead) begin
        if (MemRead == 1)
            ReadData <= memory[Address[31:2]];    //memory read
    else
        ReadData <= 32'h00000000;
    end 
    
		  
endmodule

